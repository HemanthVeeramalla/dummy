fork is cpy of repository......
